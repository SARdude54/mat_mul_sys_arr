`timescale 1ps/1ps

// Simple register implementation
// Out becomes in every clock cycle
module delay (
	input CLK,
	input [7:0] a_in,
	output logic [7:0] a_out
	);
	
	always @(posedge CLK)
		a_out <= a_in;
	
endmodule

// Module to feed values into systolic array
// Every nth row and nth col needs n delay blocks
// (n starts at 0)
module feed #(parameter M=3) (
	input CLK,
	input logic [7:0] a_in[0:(M-1)],
	output logic [7:0] a_out[0:(M-1)]
	);
	
	// Generate delay blocks here
	genvar i, j;
	generate
		for (i = 0; i < M; i++)
		begin
			// Connections between delay blocks
			logic [7:0] conn[0:i];

			// Assign input and outputs of feed module
			assign conn[0] = a_in[i];
			assign a_out[i] = conn[i];

			for (j = 0; j < i; j++)
			begin
				delay d(
					.CLK(CLK),
					.a_in(conn[j]),
					.a_out(conn[j + 1])
					);		
			end
		
		end

	endgenerate

endmodule
